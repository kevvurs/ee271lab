library verilog;
use verilog.vl_types.all;
entity discounted_testbench is
end discounted_testbench;
