library verilog;
use verilog.vl_types.all;
entity bitcompare_testbench is
end bitcompare_testbench;
