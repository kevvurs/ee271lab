library verilog;
use verilog.vl_types.all;
entity stolen_testbench is
end stolen_testbench;
