library verilog;
use verilog.vl_types.all;
entity register_testbench is
end register_testbench;
