library verilog;
use verilog.vl_types.all;
entity storeDisplay_testbench is
end storeDisplay_testbench;
