library verilog;
use verilog.vl_types.all;
entity digit_scan_testbench is
end digit_scan_testbench;
