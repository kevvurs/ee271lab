library verilog;
use verilog.vl_types.all;
entity digitDisplay_testbench is
end digitDisplay_testbench;
