library verilog;
use verilog.vl_types.all;
entity numHex_testbench is
end numHex_testbench;
